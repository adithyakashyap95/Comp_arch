// ex stage
