module func_si_forward ();

$display ("\n..............Instruction Counts...............")

$display ("\nTotal number of instructions: %d", );
$display ("Arithmetic instructions: %d",);
$display ("Logical instructions: %d",);
$display ("Memory access instructions: %d",);
$display ("Control transfer instructions: %d",);

$display ("\n\n..............Final Register State..............");

$display ("\nProgram counter: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );
$display ("R1: %d", );

$display ("\n\n..........Final memory state...........");

$display ("\nAddress: %d, Contents: %d", );
$display ("Address: %d, Contents: %d", );
$display ("Address: %d, Contents: %d", );


$display ("\n\n..........Timing Simulator..........");

$display ("\nTotal number of clock cycles: %d", );
$display ("\nProgram Halted");
