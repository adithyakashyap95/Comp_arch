// ID stage

