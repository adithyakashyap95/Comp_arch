
$display ("\n..............Instruction Counts...............")

$display ("\nTotal number of instructions: %d", );
$display ("Arithmetic instructions: %d",);
$display ("Logical instructions: %d",);
$display ("Memory access instructions: %d",);
$display ("Control transfer instructions: %d",);

$display ("\n\n..............Final Register State..............");

$display ("\nProgram counter: %d", );
$display ("R1: %d", );
$display ("R2: %d", );
$display ("R3: %d", );
$display ("R4: %d", );
$display ("R5: %d", );
$display ("R6: %d", );
$display ("R7: %d", );
$display ("R8: %d", );
$display ("R9: %d", );
$display ("R10: %d", );
$display ("R11: %d", );
$display ("R12: %d", );

$display ("\n\n..........Final memory state...........");

$display ("\nAddress: %d, Contents: %d", );
$display ("Address: %d, Contents: %d", );
$display ("Address: %d, Contents: %d", );


$display ("\n\n..........Timing Simulator..........");

$display ("\nTotal number of clock cycles: %d", );
$display ("\nProgram Halted");
