// wb stage

`include "../rtl/struct.sv"
