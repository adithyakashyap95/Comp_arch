// SV main.sv
