// ID stage

`include "../rtl/struct.sv"

