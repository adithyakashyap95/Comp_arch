// wb stage
