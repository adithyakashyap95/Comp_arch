// DATA Foreward

`include "../rtl/struct.sv"

