// Instruction fetch stage

`include "../rtl/struct.sv"
