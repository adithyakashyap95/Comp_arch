// SV main.sv

`include "../rtl/struct.sv"
