// tb .sv
