// tb .sv

`include "../rtl/struct.sv"
