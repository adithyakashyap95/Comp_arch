// mem stage
