// data hazard

`include "../rtl/struct.sv"
