// Instruction fetch stage
