// DATA Foreward
