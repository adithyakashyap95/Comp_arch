// ex stage

`include "../rtl/struct.sv"
