// ID stage

`include "../rtl/struct.sv"

// USE STRUCTURES as in struct.sv

