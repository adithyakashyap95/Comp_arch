// data hazard
